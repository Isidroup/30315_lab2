library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity lab2 is
    port (

    );
end entity lab2;

architecture RTL of lab2 is


begin


end architecture;
