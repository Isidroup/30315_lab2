-- ==============================================================
--  Lab 2 - VHDL Template
--  Descripci�n: Esqueleto de la entidad y arquitectura.
--  TODO: Completar descripci�n funcional del dise�o.
-- ==============================================================

-- TODO: A�adir librer�as necesarias.

entity lab2 is
    port (
        -- TODO: A�adir puertos de entrada/salida (se�ales, tipos, anchos).

    );
end entity lab2;

architecture RTL of lab2 is

    -- ==========================================================
    --  Declaraciones internas
    -- ==========================================================
    -- TODO: Declarar componentes .
    -- TODO: Declarar se�ales internas.
    -- TODO: Declarar constantes y tipos.

begin

    -- ==========================================================
    --  Instancias
    -- ==========================================================
    -- TODO: Instanciar subm�dulos/componentes.

    -- ==========================================================
    --  L�gica combinacional
    -- ==========================================================
    -- TODO: Implementar el modelo con bloques combinacionales.

end architecture;

