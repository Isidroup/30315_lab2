-- ==============================================================
--  Lab 2 - VHDL Template
--  Descripción: Esqueleto de la entidad y arquitectura.
--  TODO: Completar descripción funcional del diseño.
-- ==============================================================

-- TODO: Añadir librerías necesarias.

entity lab2 is
    port (
        -- TODO: Añadir puertos de entrada/salida (señales, tipos, anchos).

    );
end entity lab2;

architecture RTL of lab2 is

    -- ==========================================================
    --  Declaraciones internas
    -- ==========================================================
    -- TODO: Declarar componentes .
    -- TODO: Declarar señales internas.
    -- TODO: Declarar constantes y tipos.

begin

    -- ==========================================================
    --  Instancias
    -- ==========================================================
    -- TODO: Instanciar submódulos/componentes.

    -- ==========================================================
    --  Lógica combinacional
    -- ==========================================================
    -- TODO: Implementar el modelo con bloques combinacionales.

end architecture;
